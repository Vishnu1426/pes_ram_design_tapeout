VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pes_ram_design_tapeout
  CLASS BLOCK ;
  FOREIGN pes_ram_design_tapeout ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1800.000 ;
  PIN addr_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 115.640 1000.000 116.240 ;
    END
  END addr_a[0]
  PIN addr_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 311.480 1000.000 312.080 ;
    END
  END addr_a[1]
  PIN addr_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 507.320 1000.000 507.920 ;
    END
  END addr_a[2]
  PIN addr_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 703.160 1000.000 703.760 ;
    END
  END addr_a[3]
  PIN addr_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 899.000 1000.000 899.600 ;
    END
  END addr_a[4]
  PIN addr_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1094.840 1000.000 1095.440 ;
    END
  END addr_a[5]
  PIN addr_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 148.280 1000.000 148.880 ;
    END
  END addr_b[0]
  PIN addr_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 344.120 1000.000 344.720 ;
    END
  END addr_b[1]
  PIN addr_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 539.960 1000.000 540.560 ;
    END
  END addr_b[2]
  PIN addr_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 735.800 1000.000 736.400 ;
    END
  END addr_b[3]
  PIN addr_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 931.640 1000.000 932.240 ;
    END
  END addr_b[4]
  PIN addr_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1127.480 1000.000 1128.080 ;
    END
  END addr_b[5]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 996.000 17.720 1000.000 18.320 ;
    END
  END clk
  PIN data_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 180.920 1000.000 181.520 ;
    END
  END data_a[0]
  PIN data_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 376.760 1000.000 377.360 ;
    END
  END data_a[1]
  PIN data_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 572.600 1000.000 573.200 ;
    END
  END data_a[2]
  PIN data_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 768.440 1000.000 769.040 ;
    END
  END data_a[3]
  PIN data_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 964.280 1000.000 964.880 ;
    END
  END data_a[4]
  PIN data_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1160.120 1000.000 1160.720 ;
    END
  END data_a[5]
  PIN data_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1290.680 1000.000 1291.280 ;
    END
  END data_a[6]
  PIN data_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1421.240 1000.000 1421.840 ;
    END
  END data_a[7]
  PIN data_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 213.560 1000.000 214.160 ;
    END
  END data_b[0]
  PIN data_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 409.400 1000.000 410.000 ;
    END
  END data_b[1]
  PIN data_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 605.240 1000.000 605.840 ;
    END
  END data_b[2]
  PIN data_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 801.080 1000.000 801.680 ;
    END
  END data_b[3]
  PIN data_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 996.920 1000.000 997.520 ;
    END
  END data_b[4]
  PIN data_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1192.760 1000.000 1193.360 ;
    END
  END data_b[5]
  PIN data_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1323.320 1000.000 1323.920 ;
    END
  END data_b[6]
  PIN data_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1453.880 1000.000 1454.480 ;
    END
  END data_b[7]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1551.800 1000.000 1552.400 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.280 4.000 1236.880 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1584.440 1000.000 1585.040 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1617.080 1000.000 1617.680 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1649.720 1000.000 1650.320 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1682.360 1000.000 1682.960 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1715.000 1000.000 1715.600 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1747.640 1000.000 1748.240 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1780.280 1000.000 1780.880 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1685.080 4.000 1685.680 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1460.680 4.000 1461.280 ;
    END
  END io_oeb[9]
  PIN q_a[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 246.200 1000.000 246.800 ;
    END
  END q_a[0]
  PIN q_a[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 442.040 1000.000 442.640 ;
    END
  END q_a[1]
  PIN q_a[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 637.880 1000.000 638.480 ;
    END
  END q_a[2]
  PIN q_a[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 833.720 1000.000 834.320 ;
    END
  END q_a[3]
  PIN q_a[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1029.560 1000.000 1030.160 ;
    END
  END q_a[4]
  PIN q_a[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1225.400 1000.000 1226.000 ;
    END
  END q_a[5]
  PIN q_a[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1355.960 1000.000 1356.560 ;
    END
  END q_a[6]
  PIN q_a[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1486.520 1000.000 1487.120 ;
    END
  END q_a[7]
  PIN q_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 278.840 1000.000 279.440 ;
    END
  END q_b[0]
  PIN q_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 474.680 1000.000 475.280 ;
    END
  END q_b[1]
  PIN q_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 670.520 1000.000 671.120 ;
    END
  END q_b[2]
  PIN q_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 866.360 1000.000 866.960 ;
    END
  END q_b[3]
  PIN q_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1062.200 1000.000 1062.800 ;
    END
  END q_b[4]
  PIN q_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1258.040 1000.000 1258.640 ;
    END
  END q_b[5]
  PIN q_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1388.600 1000.000 1389.200 ;
    END
  END q_b[6]
  PIN q_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 1519.160 1000.000 1519.760 ;
    END
  END q_b[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1787.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1787.280 ;
    END
  END vssd1
  PIN we_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 50.360 1000.000 50.960 ;
    END
  END we_a
  PIN we_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 83.000 1000.000 83.600 ;
    END
  END we_b
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 1787.125 ;
      LAYER met1 ;
        RECT 4.670 10.640 999.970 1787.280 ;
      LAYER met2 ;
        RECT 4.690 10.695 999.950 1787.225 ;
      LAYER met3 ;
        RECT 4.000 1781.280 999.975 1787.205 ;
        RECT 4.000 1779.880 995.600 1781.280 ;
        RECT 4.000 1748.640 999.975 1779.880 ;
        RECT 4.000 1747.240 995.600 1748.640 ;
        RECT 4.000 1716.000 999.975 1747.240 ;
        RECT 4.000 1714.600 995.600 1716.000 ;
        RECT 4.000 1686.080 999.975 1714.600 ;
        RECT 4.400 1684.680 999.975 1686.080 ;
        RECT 4.000 1683.360 999.975 1684.680 ;
        RECT 4.000 1681.960 995.600 1683.360 ;
        RECT 4.000 1650.720 999.975 1681.960 ;
        RECT 4.000 1649.320 995.600 1650.720 ;
        RECT 4.000 1618.080 999.975 1649.320 ;
        RECT 4.000 1616.680 995.600 1618.080 ;
        RECT 4.000 1585.440 999.975 1616.680 ;
        RECT 4.000 1584.040 995.600 1585.440 ;
        RECT 4.000 1552.800 999.975 1584.040 ;
        RECT 4.000 1551.400 995.600 1552.800 ;
        RECT 4.000 1520.160 999.975 1551.400 ;
        RECT 4.000 1518.760 995.600 1520.160 ;
        RECT 4.000 1487.520 999.975 1518.760 ;
        RECT 4.000 1486.120 995.600 1487.520 ;
        RECT 4.000 1461.680 999.975 1486.120 ;
        RECT 4.400 1460.280 999.975 1461.680 ;
        RECT 4.000 1454.880 999.975 1460.280 ;
        RECT 4.000 1453.480 995.600 1454.880 ;
        RECT 4.000 1422.240 999.975 1453.480 ;
        RECT 4.000 1420.840 995.600 1422.240 ;
        RECT 4.000 1389.600 999.975 1420.840 ;
        RECT 4.000 1388.200 995.600 1389.600 ;
        RECT 4.000 1356.960 999.975 1388.200 ;
        RECT 4.000 1355.560 995.600 1356.960 ;
        RECT 4.000 1324.320 999.975 1355.560 ;
        RECT 4.000 1322.920 995.600 1324.320 ;
        RECT 4.000 1291.680 999.975 1322.920 ;
        RECT 4.000 1290.280 995.600 1291.680 ;
        RECT 4.000 1259.040 999.975 1290.280 ;
        RECT 4.000 1257.640 995.600 1259.040 ;
        RECT 4.000 1237.280 999.975 1257.640 ;
        RECT 4.400 1235.880 999.975 1237.280 ;
        RECT 4.000 1226.400 999.975 1235.880 ;
        RECT 4.000 1225.000 995.600 1226.400 ;
        RECT 4.000 1193.760 999.975 1225.000 ;
        RECT 4.000 1192.360 995.600 1193.760 ;
        RECT 4.000 1161.120 999.975 1192.360 ;
        RECT 4.000 1159.720 995.600 1161.120 ;
        RECT 4.000 1128.480 999.975 1159.720 ;
        RECT 4.000 1127.080 995.600 1128.480 ;
        RECT 4.000 1095.840 999.975 1127.080 ;
        RECT 4.000 1094.440 995.600 1095.840 ;
        RECT 4.000 1063.200 999.975 1094.440 ;
        RECT 4.000 1061.800 995.600 1063.200 ;
        RECT 4.000 1030.560 999.975 1061.800 ;
        RECT 4.000 1029.160 995.600 1030.560 ;
        RECT 4.000 1012.880 999.975 1029.160 ;
        RECT 4.400 1011.480 999.975 1012.880 ;
        RECT 4.000 997.920 999.975 1011.480 ;
        RECT 4.000 996.520 995.600 997.920 ;
        RECT 4.000 965.280 999.975 996.520 ;
        RECT 4.000 963.880 995.600 965.280 ;
        RECT 4.000 932.640 999.975 963.880 ;
        RECT 4.000 931.240 995.600 932.640 ;
        RECT 4.000 900.000 999.975 931.240 ;
        RECT 4.000 898.600 995.600 900.000 ;
        RECT 4.000 867.360 999.975 898.600 ;
        RECT 4.000 865.960 995.600 867.360 ;
        RECT 4.000 834.720 999.975 865.960 ;
        RECT 4.000 833.320 995.600 834.720 ;
        RECT 4.000 802.080 999.975 833.320 ;
        RECT 4.000 800.680 995.600 802.080 ;
        RECT 4.000 788.480 999.975 800.680 ;
        RECT 4.400 787.080 999.975 788.480 ;
        RECT 4.000 769.440 999.975 787.080 ;
        RECT 4.000 768.040 995.600 769.440 ;
        RECT 4.000 736.800 999.975 768.040 ;
        RECT 4.000 735.400 995.600 736.800 ;
        RECT 4.000 704.160 999.975 735.400 ;
        RECT 4.000 702.760 995.600 704.160 ;
        RECT 4.000 671.520 999.975 702.760 ;
        RECT 4.000 670.120 995.600 671.520 ;
        RECT 4.000 638.880 999.975 670.120 ;
        RECT 4.000 637.480 995.600 638.880 ;
        RECT 4.000 606.240 999.975 637.480 ;
        RECT 4.000 604.840 995.600 606.240 ;
        RECT 4.000 573.600 999.975 604.840 ;
        RECT 4.000 572.200 995.600 573.600 ;
        RECT 4.000 564.080 999.975 572.200 ;
        RECT 4.400 562.680 999.975 564.080 ;
        RECT 4.000 540.960 999.975 562.680 ;
        RECT 4.000 539.560 995.600 540.960 ;
        RECT 4.000 508.320 999.975 539.560 ;
        RECT 4.000 506.920 995.600 508.320 ;
        RECT 4.000 475.680 999.975 506.920 ;
        RECT 4.000 474.280 995.600 475.680 ;
        RECT 4.000 443.040 999.975 474.280 ;
        RECT 4.000 441.640 995.600 443.040 ;
        RECT 4.000 410.400 999.975 441.640 ;
        RECT 4.000 409.000 995.600 410.400 ;
        RECT 4.000 377.760 999.975 409.000 ;
        RECT 4.000 376.360 995.600 377.760 ;
        RECT 4.000 345.120 999.975 376.360 ;
        RECT 4.000 343.720 995.600 345.120 ;
        RECT 4.000 339.680 999.975 343.720 ;
        RECT 4.400 338.280 999.975 339.680 ;
        RECT 4.000 312.480 999.975 338.280 ;
        RECT 4.000 311.080 995.600 312.480 ;
        RECT 4.000 279.840 999.975 311.080 ;
        RECT 4.000 278.440 995.600 279.840 ;
        RECT 4.000 247.200 999.975 278.440 ;
        RECT 4.000 245.800 995.600 247.200 ;
        RECT 4.000 214.560 999.975 245.800 ;
        RECT 4.000 213.160 995.600 214.560 ;
        RECT 4.000 181.920 999.975 213.160 ;
        RECT 4.000 180.520 995.600 181.920 ;
        RECT 4.000 149.280 999.975 180.520 ;
        RECT 4.000 147.880 995.600 149.280 ;
        RECT 4.000 116.640 999.975 147.880 ;
        RECT 4.000 115.280 995.600 116.640 ;
        RECT 4.400 115.240 995.600 115.280 ;
        RECT 4.400 113.880 999.975 115.240 ;
        RECT 4.000 84.000 999.975 113.880 ;
        RECT 4.000 82.600 995.600 84.000 ;
        RECT 4.000 51.360 999.975 82.600 ;
        RECT 4.000 49.960 995.600 51.360 ;
        RECT 4.000 18.720 999.975 49.960 ;
        RECT 4.000 17.320 995.600 18.720 ;
        RECT 4.000 10.715 999.975 17.320 ;
      LAYER met4 ;
        RECT 854.975 17.855 865.440 1054.505 ;
        RECT 867.840 17.855 942.240 1054.505 ;
        RECT 944.640 17.855 998.825 1054.505 ;
  END
END pes_ram_design_tapeout
END LIBRARY

