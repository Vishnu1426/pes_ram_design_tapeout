magic
tech sky130A
magscale 1 2
timestamp 1700941454
<< obsli1 >>
rect 1104 2159 198812 357425
<< obsm1 >>
rect 934 2128 199994 357456
<< obsm2 >>
rect 938 2139 199990 357445
<< metal3 >>
rect 199200 356056 200000 356176
rect 199200 349528 200000 349648
rect 199200 343000 200000 343120
rect 0 337016 800 337136
rect 199200 336472 200000 336592
rect 199200 329944 200000 330064
rect 199200 323416 200000 323536
rect 199200 316888 200000 317008
rect 199200 310360 200000 310480
rect 199200 303832 200000 303952
rect 199200 297304 200000 297424
rect 0 292136 800 292256
rect 199200 290776 200000 290896
rect 199200 284248 200000 284368
rect 199200 277720 200000 277840
rect 199200 271192 200000 271312
rect 199200 264664 200000 264784
rect 199200 258136 200000 258256
rect 199200 251608 200000 251728
rect 0 247256 800 247376
rect 199200 245080 200000 245200
rect 199200 238552 200000 238672
rect 199200 232024 200000 232144
rect 199200 225496 200000 225616
rect 199200 218968 200000 219088
rect 199200 212440 200000 212560
rect 199200 205912 200000 206032
rect 0 202376 800 202496
rect 199200 199384 200000 199504
rect 199200 192856 200000 192976
rect 199200 186328 200000 186448
rect 199200 179800 200000 179920
rect 199200 173272 200000 173392
rect 199200 166744 200000 166864
rect 199200 160216 200000 160336
rect 0 157496 800 157616
rect 199200 153688 200000 153808
rect 199200 147160 200000 147280
rect 199200 140632 200000 140752
rect 199200 134104 200000 134224
rect 199200 127576 200000 127696
rect 199200 121048 200000 121168
rect 199200 114520 200000 114640
rect 0 112616 800 112736
rect 199200 107992 200000 108112
rect 199200 101464 200000 101584
rect 199200 94936 200000 95056
rect 199200 88408 200000 88528
rect 199200 81880 200000 82000
rect 199200 75352 200000 75472
rect 199200 68824 200000 68944
rect 0 67736 800 67856
rect 199200 62296 200000 62416
rect 199200 55768 200000 55888
rect 199200 49240 200000 49360
rect 199200 42712 200000 42832
rect 199200 36184 200000 36304
rect 199200 29656 200000 29776
rect 199200 23128 200000 23248
rect 0 22856 800 22976
rect 199200 16600 200000 16720
rect 199200 10072 200000 10192
rect 199200 3544 200000 3664
<< obsm3 >>
rect 800 356256 199995 357441
rect 800 355976 199120 356256
rect 800 349728 199995 355976
rect 800 349448 199120 349728
rect 800 343200 199995 349448
rect 800 342920 199120 343200
rect 800 337216 199995 342920
rect 880 336936 199995 337216
rect 800 336672 199995 336936
rect 800 336392 199120 336672
rect 800 330144 199995 336392
rect 800 329864 199120 330144
rect 800 323616 199995 329864
rect 800 323336 199120 323616
rect 800 317088 199995 323336
rect 800 316808 199120 317088
rect 800 310560 199995 316808
rect 800 310280 199120 310560
rect 800 304032 199995 310280
rect 800 303752 199120 304032
rect 800 297504 199995 303752
rect 800 297224 199120 297504
rect 800 292336 199995 297224
rect 880 292056 199995 292336
rect 800 290976 199995 292056
rect 800 290696 199120 290976
rect 800 284448 199995 290696
rect 800 284168 199120 284448
rect 800 277920 199995 284168
rect 800 277640 199120 277920
rect 800 271392 199995 277640
rect 800 271112 199120 271392
rect 800 264864 199995 271112
rect 800 264584 199120 264864
rect 800 258336 199995 264584
rect 800 258056 199120 258336
rect 800 251808 199995 258056
rect 800 251528 199120 251808
rect 800 247456 199995 251528
rect 880 247176 199995 247456
rect 800 245280 199995 247176
rect 800 245000 199120 245280
rect 800 238752 199995 245000
rect 800 238472 199120 238752
rect 800 232224 199995 238472
rect 800 231944 199120 232224
rect 800 225696 199995 231944
rect 800 225416 199120 225696
rect 800 219168 199995 225416
rect 800 218888 199120 219168
rect 800 212640 199995 218888
rect 800 212360 199120 212640
rect 800 206112 199995 212360
rect 800 205832 199120 206112
rect 800 202576 199995 205832
rect 880 202296 199995 202576
rect 800 199584 199995 202296
rect 800 199304 199120 199584
rect 800 193056 199995 199304
rect 800 192776 199120 193056
rect 800 186528 199995 192776
rect 800 186248 199120 186528
rect 800 180000 199995 186248
rect 800 179720 199120 180000
rect 800 173472 199995 179720
rect 800 173192 199120 173472
rect 800 166944 199995 173192
rect 800 166664 199120 166944
rect 800 160416 199995 166664
rect 800 160136 199120 160416
rect 800 157696 199995 160136
rect 880 157416 199995 157696
rect 800 153888 199995 157416
rect 800 153608 199120 153888
rect 800 147360 199995 153608
rect 800 147080 199120 147360
rect 800 140832 199995 147080
rect 800 140552 199120 140832
rect 800 134304 199995 140552
rect 800 134024 199120 134304
rect 800 127776 199995 134024
rect 800 127496 199120 127776
rect 800 121248 199995 127496
rect 800 120968 199120 121248
rect 800 114720 199995 120968
rect 800 114440 199120 114720
rect 800 112816 199995 114440
rect 880 112536 199995 112816
rect 800 108192 199995 112536
rect 800 107912 199120 108192
rect 800 101664 199995 107912
rect 800 101384 199120 101664
rect 800 95136 199995 101384
rect 800 94856 199120 95136
rect 800 88608 199995 94856
rect 800 88328 199120 88608
rect 800 82080 199995 88328
rect 800 81800 199120 82080
rect 800 75552 199995 81800
rect 800 75272 199120 75552
rect 800 69024 199995 75272
rect 800 68744 199120 69024
rect 800 67936 199995 68744
rect 880 67656 199995 67936
rect 800 62496 199995 67656
rect 800 62216 199120 62496
rect 800 55968 199995 62216
rect 800 55688 199120 55968
rect 800 49440 199995 55688
rect 800 49160 199120 49440
rect 800 42912 199995 49160
rect 800 42632 199120 42912
rect 800 36384 199995 42632
rect 800 36104 199120 36384
rect 800 29856 199995 36104
rect 800 29576 199120 29856
rect 800 23328 199995 29576
rect 800 23056 199120 23328
rect 880 23048 199120 23056
rect 880 22776 199995 23048
rect 800 16800 199995 22776
rect 800 16520 199120 16800
rect 800 10272 199995 16520
rect 800 9992 199120 10272
rect 800 3744 199995 9992
rect 800 3464 199120 3744
rect 800 2143 199995 3464
<< metal4 >>
rect 4208 2128 4528 357456
rect 19568 2128 19888 357456
rect 34928 2128 35248 357456
rect 50288 2128 50608 357456
rect 65648 2128 65968 357456
rect 81008 2128 81328 357456
rect 96368 2128 96688 357456
rect 111728 2128 112048 357456
rect 127088 2128 127408 357456
rect 142448 2128 142768 357456
rect 157808 2128 158128 357456
rect 173168 2128 173488 357456
rect 188528 2128 188848 357456
<< obsm4 >>
rect 170995 3571 173088 210901
rect 173568 3571 188448 210901
rect 188928 3571 199765 210901
<< labels >>
rlabel metal3 s 199200 23128 200000 23248 6 addr_a[0]
port 1 nsew signal input
rlabel metal3 s 199200 62296 200000 62416 6 addr_a[1]
port 2 nsew signal input
rlabel metal3 s 199200 101464 200000 101584 6 addr_a[2]
port 3 nsew signal input
rlabel metal3 s 199200 140632 200000 140752 6 addr_a[3]
port 4 nsew signal input
rlabel metal3 s 199200 179800 200000 179920 6 addr_a[4]
port 5 nsew signal input
rlabel metal3 s 199200 218968 200000 219088 6 addr_a[5]
port 6 nsew signal input
rlabel metal3 s 199200 29656 200000 29776 6 addr_b[0]
port 7 nsew signal input
rlabel metal3 s 199200 68824 200000 68944 6 addr_b[1]
port 8 nsew signal input
rlabel metal3 s 199200 107992 200000 108112 6 addr_b[2]
port 9 nsew signal input
rlabel metal3 s 199200 147160 200000 147280 6 addr_b[3]
port 10 nsew signal input
rlabel metal3 s 199200 186328 200000 186448 6 addr_b[4]
port 11 nsew signal input
rlabel metal3 s 199200 225496 200000 225616 6 addr_b[5]
port 12 nsew signal input
rlabel metal3 s 199200 3544 200000 3664 6 clk
port 13 nsew signal input
rlabel metal3 s 199200 36184 200000 36304 6 data_a[0]
port 14 nsew signal input
rlabel metal3 s 199200 75352 200000 75472 6 data_a[1]
port 15 nsew signal input
rlabel metal3 s 199200 114520 200000 114640 6 data_a[2]
port 16 nsew signal input
rlabel metal3 s 199200 153688 200000 153808 6 data_a[3]
port 17 nsew signal input
rlabel metal3 s 199200 192856 200000 192976 6 data_a[4]
port 18 nsew signal input
rlabel metal3 s 199200 232024 200000 232144 6 data_a[5]
port 19 nsew signal input
rlabel metal3 s 199200 258136 200000 258256 6 data_a[6]
port 20 nsew signal input
rlabel metal3 s 199200 284248 200000 284368 6 data_a[7]
port 21 nsew signal input
rlabel metal3 s 199200 42712 200000 42832 6 data_b[0]
port 22 nsew signal input
rlabel metal3 s 199200 81880 200000 82000 6 data_b[1]
port 23 nsew signal input
rlabel metal3 s 199200 121048 200000 121168 6 data_b[2]
port 24 nsew signal input
rlabel metal3 s 199200 160216 200000 160336 6 data_b[3]
port 25 nsew signal input
rlabel metal3 s 199200 199384 200000 199504 6 data_b[4]
port 26 nsew signal input
rlabel metal3 s 199200 238552 200000 238672 6 data_b[5]
port 27 nsew signal input
rlabel metal3 s 199200 264664 200000 264784 6 data_b[6]
port 28 nsew signal input
rlabel metal3 s 199200 290776 200000 290896 6 data_b[7]
port 29 nsew signal input
rlabel metal3 s 199200 310360 200000 310480 6 io_oeb[0]
port 30 nsew signal output
rlabel metal3 s 0 247256 800 247376 6 io_oeb[10]
port 31 nsew signal output
rlabel metal3 s 0 202376 800 202496 6 io_oeb[11]
port 32 nsew signal output
rlabel metal3 s 0 157496 800 157616 6 io_oeb[12]
port 33 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 io_oeb[13]
port 34 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 io_oeb[14]
port 35 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 io_oeb[15]
port 36 nsew signal output
rlabel metal3 s 199200 316888 200000 317008 6 io_oeb[1]
port 37 nsew signal output
rlabel metal3 s 199200 323416 200000 323536 6 io_oeb[2]
port 38 nsew signal output
rlabel metal3 s 199200 329944 200000 330064 6 io_oeb[3]
port 39 nsew signal output
rlabel metal3 s 199200 336472 200000 336592 6 io_oeb[4]
port 40 nsew signal output
rlabel metal3 s 199200 343000 200000 343120 6 io_oeb[5]
port 41 nsew signal output
rlabel metal3 s 199200 349528 200000 349648 6 io_oeb[6]
port 42 nsew signal output
rlabel metal3 s 199200 356056 200000 356176 6 io_oeb[7]
port 43 nsew signal output
rlabel metal3 s 0 337016 800 337136 6 io_oeb[8]
port 44 nsew signal output
rlabel metal3 s 0 292136 800 292256 6 io_oeb[9]
port 45 nsew signal output
rlabel metal3 s 199200 49240 200000 49360 6 q_a[0]
port 46 nsew signal output
rlabel metal3 s 199200 88408 200000 88528 6 q_a[1]
port 47 nsew signal output
rlabel metal3 s 199200 127576 200000 127696 6 q_a[2]
port 48 nsew signal output
rlabel metal3 s 199200 166744 200000 166864 6 q_a[3]
port 49 nsew signal output
rlabel metal3 s 199200 205912 200000 206032 6 q_a[4]
port 50 nsew signal output
rlabel metal3 s 199200 245080 200000 245200 6 q_a[5]
port 51 nsew signal output
rlabel metal3 s 199200 271192 200000 271312 6 q_a[6]
port 52 nsew signal output
rlabel metal3 s 199200 297304 200000 297424 6 q_a[7]
port 53 nsew signal output
rlabel metal3 s 199200 55768 200000 55888 6 q_b[0]
port 54 nsew signal output
rlabel metal3 s 199200 94936 200000 95056 6 q_b[1]
port 55 nsew signal output
rlabel metal3 s 199200 134104 200000 134224 6 q_b[2]
port 56 nsew signal output
rlabel metal3 s 199200 173272 200000 173392 6 q_b[3]
port 57 nsew signal output
rlabel metal3 s 199200 212440 200000 212560 6 q_b[4]
port 58 nsew signal output
rlabel metal3 s 199200 251608 200000 251728 6 q_b[5]
port 59 nsew signal output
rlabel metal3 s 199200 277720 200000 277840 6 q_b[6]
port 60 nsew signal output
rlabel metal3 s 199200 303832 200000 303952 6 q_b[7]
port 61 nsew signal output
rlabel metal4 s 4208 2128 4528 357456 6 vccd1
port 62 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 357456 6 vccd1
port 62 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 357456 6 vccd1
port 62 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 357456 6 vccd1
port 62 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 357456 6 vccd1
port 62 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 357456 6 vccd1
port 62 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 357456 6 vccd1
port 62 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 357456 6 vssd1
port 63 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 357456 6 vssd1
port 63 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 357456 6 vssd1
port 63 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 357456 6 vssd1
port 63 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 357456 6 vssd1
port 63 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 357456 6 vssd1
port 63 nsew ground bidirectional
rlabel metal3 s 199200 10072 200000 10192 6 we_a
port 64 nsew signal input
rlabel metal3 s 199200 16600 200000 16720 6 we_b
port 65 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 200000 360000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 30725812
string GDS_FILE /home/vishnu/pes_ram_design_tapeout/openlane/pes_ram_design_tapeout/runs/23_11_26_01_03/results/signoff/pes_ram_design_tapeout.magic.gds
string GDS_START 555344
<< end >>

